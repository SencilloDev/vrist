module vrist 

